module RF_256_64 ( CLK, CEB, WEB, A, D, BWEB, Q );

parameter numWord = 256;
parameter numRow = 64;
parameter numCM = 4;
parameter numBit = 64;
parameter numWordAddr = 8;
parameter numRowAddr = 6;
parameter numCMAddr = 2;
	
// this is a proprietary model and cannot be shared openly. we make the parameters available above for reference.

endmodule
`endcelldefine


