`timescale 1ns / 1ps

/************************************************************************************************
    1. Design Name:             tb_kem_dec_cca
    2. Preparation Date:        June 02, 2021
    3. Initial designed by:     Malik Imran and Samuel Pagliarini (Tallinn University of Technology, Estonia)              
    
    Note! The codes are for academic research use only and does not come with any support or any responsibility. 
****************************************************************************************************/

module tb_kem_dec_cca;

	// Inputs to the core
	reg clk1;
	reg clk2;
	reg rst;
	reg addr;
	reg din;
	reg addr_ready;
	reg LAD1;
	reg LAD2;
	reg we;
    reg CONT;
    reg start;	
    reg crypto_op_1;
    reg crypto_op_2;
    reg crypto_op_3;
    	
	// Outputs from the core
	wire dout;
	wire done;
    
	// Registers declaration to hold the test values and signals (i.e., i and count) to drive loops (i.e., for) to read values
	reg [10:0] i;
	reg [9:0] j, count;	
	reg [63:0] set_memory;
	reg [63:0] cpa_secret[47:0];	// 3 secret polynomials where each coeff is in signed magnitude and occupies 4 bits
	reg [63:0] pk[123:0];			// 120 words are for CPA pk and the next 4 words are seed_A
	reg [63:0] hash_pk[3:0];		// 4 words are for hash(pk)	
	reg [63:0] pseudo_random[3:0]; 	// If decapsulation fails, this pseudo_random string is output
	reg [63:0] ct[135:0];			// 960 + 128 bytes
	reg [63:0] last_data_on_last_memory_address;
	reg [6:0]  counter_to_read_64_bit_segment;
	
	// Instantiate the Unit Under Test (UUT)	
	wrapper_top uut (
		.clk1(clk1),
		.clk2(clk2), 
		.rst(rst),
		.addr(addr), 
		.din(din), 
		.addr_ready(addr_ready),
		.LAD1(LAD1),
	    .LAD2(LAD2),
	    .we(we),
	    .CONT(CONT),
	    .start(start),
	    .crypto_op_1(crypto_op_1),
	    .crypto_op_2(crypto_op_2), 
	    .crypto_op_3(crypto_op_3),
		.dout(dout),
		.done(done)     		
	);

	initial begin
		// Initialize Inputs
		clk1 = 0;
		clk2 = 0;
		rst = 1;
		addr = 0;
		din = 0;
		addr_ready = 0;
		LAD1 = 0;
		LAD2 = 0;
		we = 0;
		CONT = 0;
		start = 0;
		crypto_op_1 = 0;
	    crypto_op_2 = 0;
	    crypto_op_3 = 0;
	    
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%%      Test vectors for the Decapsulation 
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/	

		cpa_secret[0] = 64'b1001001110011010000100000001100100000001001010100000000010010001;//h939a1019012a0091;
		cpa_secret[1] = 64'b000110010000000010010010001000010000001000010011100110111010;//h1900922102139ba;
		cpa_secret[2] = 64'b1011101000001011101000000001100100001001000000010000110000001010;//hba0ba01909010c0a;
		cpa_secret[3] = 64'b0010000100010000100110010000000000011010100110010000100110011001;//h211099001a990999;
		cpa_secret[4] = 64'b1001100100010001001100010001000100000000000010010010000100010000;//'h9911311100092110;
		cpa_secret[5] = 64'b000110101010000010100001100100011010000010010001100100011011;//h1aa0a191a09191b;
		cpa_secret[6] = 64'b101010110001000110010000000100001001100100010001000000000000;//hab1190109911000;
		cpa_secret[7] = 64'b101010111001000100010001000000110001000010100010000010100011;//hab91110310a20a3;
		cpa_secret[8] = 64'b0011101000010100000010010010100100000001101010011001000100001010;//h3a14092901a9910a;
		cpa_secret[9] = 64'b1001001000001001000010011010000000001001000000110010000100101001;//h920909a009032129;
		cpa_secret[10] = 64'b101010011010000100100000001000000010000010111001101000010001;//ha9a1202020b9a11;
		cpa_secret[11] = 64'b1001001000000000000000010001000100011010000000001010001110010000;//h920001111a00a390;
		cpa_secret[12] = 64'b100110011010000000001010101100010000000110010001000000011001;//h99a00ab10191019;
		cpa_secret[13] = 64'b100100011010000000101010000110101010001000010001100100010001;//h91a02a1aa211911;
		cpa_secret[14] = 64'b0001100110010000100100000000000100011010001010101001000110011001;//h199090011a2a9199;
		cpa_secret[15] = 64'b0001100100000000100100010001001000011001001000010000100100010010;//h1900911219210912;
		cpa_secret[16] = 64'b0001101000000001000000011001001100010000000010010001000000001001;//h1a01019310091009;
		cpa_secret[17] = 64'b1011101000110001000000000001100100011011100100101001101000010001;//hba3100191b929a11;
		cpa_secret[18] = 64'b0001000000100001000000000000000000010000101000001001000000000000;//h1021000010a09000;
		cpa_secret[19] = 64'b1010000000001010000000100010000100010010101010100010100100001011;//ha00a022112aa290b;
		cpa_secret[20] = 64'b1001100100100010100100100001000010100001000100010010000100010001;//h99229210a1112111;
		cpa_secret[21] = 64'b100110010000000100000001000000000000000110100000000000111001;//h9901010001a0039;
		cpa_secret[22] = 64'b0010001010010000101010010010101000001001100100010001;//h2290a92a09911;
		cpa_secret[23] = 64'b0001000110010001000100100000000010010000000100000000100100000000;//h1191120090100900;
		cpa_secret[24] = 64'b1010000000111001000000010000000000101001100100110001100100110000;//ha039010029931930;
		cpa_secret[25] = 64'b0001000110010000000000001001000100010010101100010010101000001010;//h1190009112b12a0a;
		cpa_secret[26] = 64'b000100011001101000010001001000000000000100111001001000101010;//h119a1120013922a;
		cpa_secret[27] = 64'b001000010001101100011010100110101001001010111001000110010000;//h211b1a9a92b9190;
		cpa_secret[28] = 64'b0001001100000001000110011001100100010000000000010001;//h1301199910011;
		cpa_secret[29] = 64'b0001000010110001000100100010000000101001000110101001001000001001;//h10b11220291a9209;
		cpa_secret[30] = 64'b0001100110010000000100010000000000100001000100000010000000000000;//h1990110021102000;
		cpa_secret[31] = 64'b1010000010010001000100101001000010101001101010010100101000100000;//ha0911290a9a94a20;
		cpa_secret[32] = 64'b000110011001100100000010000010101010101000001001001000001010;//h1999020aaa0920a;
		cpa_secret[33] = 64'b1001100110010001000100100010101100011010000000110010;//h9991122b1a032;
		cpa_secret[34] = 64'b0001000100010000000110110010000010011010101000010001000100000000;//h11101b209aa11100;
		cpa_secret[35] = 64'b0001100100010001101000000010100110101001100100101011000110011001;//h1911a029a992b199;
		cpa_secret[36] = 64'b0001101100011010000000010000000110010000000000010010000110011100;//h1b1a01019001219c;
		cpa_secret[37] = 64'b0001000010010000101000100000101010010010100100011010100100000001;//h1090a20a9291a901;
		cpa_secret[38] = 64'b101010010000100110010000000100010001000110101001001011000001;//ha909901111a92c1;
		cpa_secret[39] = 64'b1001101000101010100100001001000010010000001010100000001100011010;//h9a2a9090902a031a;
		cpa_secret[40] = 64'b1010100100000000100110010001000110110000100110110000101000101001;//ha9009911b09b0a29;
		cpa_secret[41] = 64'b1001000000000000000100001001000110011001101010100001101100011010;//h9000109199aa1b1a;
		cpa_secret[42] = 64'b1010000010011010000010100001000100010001001110010001001000010000;//ha09a0a1111391210;
		cpa_secret[43] = 64'b0001000100001001000000010001000110010001000000011001100110011010;//h110901119101999a;
		cpa_secret[44] = 64'b1010000000010001000000010001101000010000001000010010100100011001;//ha011011a10212919;
		cpa_secret[45] = 64'b001000000001000100010001000000000001100100110010000000010010;//h201111001932012;
		cpa_secret[46] = 64'b1010100110101010100110011010000000010000100100010010101000011001;//ha9aa99a010912a19;
		cpa_secret[47] = 64'b0010000110101001000000011001100100011001101000001010100100000010;//h21a9019919a0a902;

        // 120+4 word pk 
		pk[0] = 64'b1101101100001100101101100111101000010111101010011010111011101011;//hdb0cb67a17a9aeeb;
		pk[1] = 64'b1010111100011001100111111001011011011111101101101110010100100001;//haf199f96dfb6e521;
		pk[2] = 64'b1010100001001100000010110000010110100011000111110000011101110011;//ha84c0b05a31f0773;
		pk[3] = 64'b1110010011100111010110100011100011111110100110110111111010010000;//he4e75a38fe9b7e90;
		pk[4] = 64'b1000001100000110001110111011111101001010101101101111000111101001;//h83063bbf4ab6f1e9;
		pk[5] = 64'b1100111000100100101001111101001101000110000100101001110101100001;//hce24a7d346129d61;
		pk[6] = 64'b0101100111011000011000100111011110110101110001001001001100101100;//h59d86277b5c4932c;
		pk[7] = 64'b1010101011101000010000100110100110001001101000101011111001000111;//haae8426989a2be47;
		pk[8] = 64'b1010001001010001101110101111111111110011101100100111101100011110;//ha251bafff3b27b1e;
		pk[9] =  64'b1100011110101000110000110011001110010001011111111101100110010110;//hc7a8c333917fd996;
		pk[10] = 64'b0010010010110101111001011000110111100011000110001111110101001101;//h24b5e58de318fd4d;
		pk[11] = 64'b1000010000000101011010001001000110000101111010000100000100001110;//h8405689185e8410e;
		pk[12] = 64'b0101001010010000110100011001110011011111010111001100011000100100;//h5290d19cdf5cc624;
		pk[13] = 64'b1000010100011111011100101111011101011010100010101111100000000010;//h851f72f75a8af802;
		pk[14] = 64'b0111110110111001001001111111100111110010011101000100000100000110;//h7db927f9f2744106;
		pk[15] = 64'b0001111110100010000111110010011001011111110011101000000101101001;//h1fa21f265fce8169;
		pk[16] = 64'b0010001110110011011110010011101110111011011101001011111011111010;//h23b3793bbb74befa;
		pk[17] = 64'b1000000110100110101001100000010110100111001000100100100010100101;//h81a6a605a72248a5;
		pk[18] = 64'b0101110010011111011110101111001111010001111011101100001001010111;//h5c9f7af3d1eec257;
		pk[19] = 64'b0011010110111010110000010110011110100110110101011010000101101001;//h35bac167a6d5a169;
		pk[20] = 64'b1011101100110111000111111101001011110001011011111011111111010100;//hbb371fd2f16fbfd4;
		pk[21] = 64'b0011101001001011111011101101110101010101100100110000111000001001;//h3a4beedd55930e09;
		pk[22] = 64'b1010011110110000101000010011100011101000110011001010100010000111;//ha7b0a138e8cca887;
		pk[23] = 64'b100010110010010010000100101101010001010001111010011111110110;//h8b2484b5147a7f6;
		pk[24] = 64'b1101110000110010101000011100110010101111011001001101001110011000;//hdc32a1ccaf64d398;
		pk[25] = 64'b0101110100100011001111000000011100010010111110110101001000001111;//h5d233c0712fb520f;
		pk[26] = 64'b0001101100001010000110110011010000000011011110110001111100101000;//h1b0a1b34037b1f28;
		pk[27] = 64'b0100000111010110110101101101110001100100111011101010011000001011;//h41d6d6dc64eea60b;
		pk[28] = 64'b0110101000101010100010000001111001000111100000100011110100111000;//h6a2a881e47823d38;
		pk[29] = 64'b1010010101010111011101010100001010101000100011101001111110010101;//ha5577542a88e9f95;
		pk[30] = 64'b1101010111010100111100000000010101100101111011101111000010100011;//hd5d4f00565eef0a3;
		pk[31] = 64'b1010100111000010111111101011011000011111000001011001100100101100;//ha9c2feb61f05992c;
		pk[32] = 64'b1010100110111000001001100110011110000011011000010111001101001110;//ha9b826678361734e;
		pk[33] = 64'b0101100011010000000110001001110110101000010110001111010000100111;//h58d0189da858f427;
		pk[34] = 64'b0101011111100001000110010010100011111011110000101001111010011111;//h57e11928fbc29e9f;
		pk[35] = 64'b0010100110001100011000100000101111101100011100101001011101101111;//h298c620bec72976f;
		pk[36] = 64'b1011101001101010101000101110110100110101111111000111110111101000;//hba6aa2ed35fc7de8;
		pk[37] = 64'b010110111010011011011100101010101001011001101101010100011101;//h5ba6dcaa966d51d;
		pk[38] = 64'b0101101100100010000010010110010011001111110011011001110001010001;//h5b220964cfcd9c51;
		pk[39] = 64'b0010110100001011110010100100001100111111000101010111011000011000;//h2d0bca433f157618;
		pk[40] = 64'b1001101101000100001110101010010110100101100101111001011011101111;//h9b443aa5a59796ef;
		pk[41] = 64'b0100111000000101001111111011110010100111111010101110000101000110;//h4e053fbca7eae146;
		pk[42] = 64'b1010000001101110000010001000110010110110001110101010100001011101;//ha06e088cb63aa85d;
		pk[43] = 64'b1011010011101001011001010010100100110010100011001010100111001001;//hb4e96529328ca9c9;
		pk[44] = 64'b0010001111000110100000110001101111000110010100100110110101000110;//h23c6831bc6526d46;
		pk[45] = 64'b1100100110110101010011001110000110001011101000101110111001000101;//hc9b54ce18ba2ee45;
		pk[46] = 64'b0111011001100000111011111111011100011110010001110100010101101111;//h7660eff71e47456f;
		pk[47] = 64'b1001100110001000101010001010011100111111110111111110001110101111;//h9988a8a73fdfe3af;
		pk[48] = 64'b1000100011011111101111111101110010111111001100100010111011000110;//h88dfbfdcbf322ec6;
		pk[49] = 64'b1010001000010000100011001000000000010011010001010110010010010111;//ha2108c8013456497;
		pk[50] = 64'b1110011010010100111010101111011100111000111110101011111100001001;//he694eaf738fabf09;
		pk[51] = 64'b1111111110101101101110001100001110011011000100110000111110101100;//hffadb8c39b130fac;
		pk[52] = 64'b0011110110111110001100000101011001110100001101101010111111000100;//h3dbe30567436afc4;
		pk[53] = 64'b1111111010011100100101110111111001110111001110000101000010100111;//hfe9c977e773850a7;
		pk[54] = 64'b1101110000011100000011100100011100011001101111011100010011000000;//hdc1c0e4719bdc4c0;
		pk[55] = 64'b0111000011111011010000101011001011011100100001100010100100101111;//h70fb42b2dc86292f;
		pk[56] = 64'b1011100100001101001110110111010100101110001100110101011001111111;//hb90d3b752e33567f;
		pk[57] = 64'b1111000111000010100001111001011100001000110000010110100010001110;//hf1c2879708c1688e;
		pk[58] = 64'b1000100101010010000111000000001010001110001111111011001111011011;//h89521c028e3fb3db;
		pk[59] = 64'b1110011001001111001001110110000101100101000011010100010011010110;//he64f2761650d44d6;
		pk[60] = 64'b0011101000111001110010011011111100000001100001100001010011111111;//h3a39c9bf018614ff;
		pk[61] = 64'b0111010010100010000100010001101011011111101010010101000000011010;//h74a2111adfa9501a;
		pk[62] = 64'b1100001011101001000100100100100111110000011010111000000001000111;//hc2e91249f06b8047;
		pk[63] = 64'b0100001111001001100011101011101011100111001101010011110000010000;//h43c98ebae7353c10;
		pk[64] = 64'b1001101010011111110101111010000010101110110110101011010000110010;//h9a9fd7a0aedab432;
		pk[65] = 64'b0100011010110001010101110000100101000101011111101010110100100001;//h46b15709457ead21;
		pk[66] = 64'b0100111101011110111001100111011101000111101001000011101110001101;//h4f5ee67747a43b8d;
		pk[67] = 64'b0011101100001101100100001100111010000000000100001011010000110100;//h3b0d90ce8010b434;
		pk[68] = 64'b0100011001010001101000100111000101101001111010110100011011001011;//h4651a27169eb46cb;
		pk[69] = 64'b1100100011100001101011000000110000011101101010010101101110111101;//hc8e1ac0c1da95bbd;
		pk[70] = 64'b0100100111100110101111001111000100010000011000100011101100110000;//h49e6bcf110623b30;
		pk[71] = 64'b1000101011001110011000010001000011101101100100101111110111001100;//h8ace6110ed92fdcc;
		pk[72] = 64'b1110001011011110111001011100100010001001111001101000111101000110;//he2dee5c889e68f46;
		pk[73] = 64'b1011001111000001100010000001101011110111010111000010110110001100;//hb3c1881af75c2d8c;
		pk[74] = 64'b110100101001100101111001101100000011100000100100001011111101;//hd29979b038242fd;
		pk[75] = 64'b0001110011001110111000000000001001011010110111000010001111101001;//h1ccee0025adc23e9;
		pk[76] = 64'b0111101000100010010010110101000001010100101011110110111001101111;//h7a224b5054af6e6f;
		pk[77] = 64'b1111010110011100011110010100101000011001001111000001100001000100;//hf59c794a193c1844;
		pk[78] = 64'b1000100010111011010100100110101001111101000000011111101101110000;//h88bb526a7d01fb70;
		pk[79] = 64'b1101111100010111101100111111110111000000011000101111100011011111;//hdf17b3fdc062f8df;
		pk[80] = 64'b10011001100110100101011101001100001110100101101111011011;//h999a574c3a5bdb;
		pk[81] = 64'b0110101010001010100001111100110110100000000001010100011100100011;//h6a8a87cda0054723;
		pk[82] = 64'b1000111000010101110010110100101100000110111010011111000100100011;//h8e15cb4b06e9f123;
		pk[83] = 64'b1110100100111100010111110111010101101000111001001101011110010010;//he93c5f7568e4d792;
		pk[84] = 64'b0110101111101001100100110000111000100100110110010010110001101101;//h6be9930e24d92c6d;
		pk[85] = 64'b1011011101001011011011110010001101000010011100111100011011101111;//hb74b6f234273c6ef;
		pk[86] = 64'b0110110110010101111100001001001010100101001101010101010011111110;//h6d95f092a53554fe;
		pk[87] = 64'b0110001100001001000111001100001010001001110110010111000011110010;//h63091cc289d970f2;
		pk[88] = 64'b1010110101000010111110111011001011001001010110101100011001011110;//had42fbb2c95ac65e;
		pk[89] = 64'b1111101110101101101010001110001110001001101001001101011010101011;//hfbada8e389a4d6ab;
		pk[90] = 64'b1011101001110010011111101001011001011110110001010011101111110001;//hba727e965ec53bf1;
		pk[91] = 64'b0101111010101101111101010000010010000101110011001100110110100101;//h5eadf50485cccda5;
		pk[92] = 64'b1011110000001100100011110101011011111111110011001000000011100001;//hbc0c8f56ffcc80e1;
		pk[93] = 64'b0100010111011011100100001101001011111110000000100011001111001111;//h45db90d2fe0233cf;
		pk[94] = 64'b1110110001000001110011110110100100010010100000011010110100010001;//hec41cf691281ad11;
		pk[95] = 64'b1111000101010100101100011001001001011011000011101010111010011100;//hf154b1925b0eae9c;
		pk[96] = 64'b1100111100101001111101100100110100111000110100101101010111000110;//hcf29f64d38d2d5c6;
		pk[97] = 64'b1101001100101111011111100101010011000000110110100000000010101010;//hd32f7e54c0da00aa;
		pk[98] = 64'b0011001110100000110101011101011111011010111000111111111001111100;//h33a0d5d7dae3fe7c;
		pk[99] =  64'b1110000001001101010100111010111011001101110011000011011111110110;//he04d53aecdcc37f6;
		pk[100] = 64'b0001011111010110100001110011110100101010100100101110011000001001;//h17d6873d2a92e609;
		pk[101] = 64'b0101111010100101010111001000100001010010010001100110011001110110;//h5ea55c8852466676;
		pk[102] = 64'b1010100101100110111011001010101110111011101010111001101010110011;//ha966ecabbbab9ab3;
		pk[103] = 64'b1100000000111101010111110100100000101101100000100111000111001101;//hc03d5f482d8271cd;
		pk[104] = 64'b0010011010111111001001010101100101101000110111011111011010100000;//h26bf255968ddf6a0;
		pk[105] = 64'b0111110011000000001011001100001001010011100010001110010000110100;//h7cc02cc25388e434;
		pk[106] = 64'b1101101100000111001111011011100101011110001111110001101010110001;//hdb073db95e3f1ab1;
		pk[107] = 64'b1110101011101000000000010011010001100011100101111000010010111001;//heae80134639784b9;
		pk[108] = 64'b001111011000011101110000110000111111101100000000011100010110;//h3d8770c3fb00716;
		pk[109] = 64'b1011001011000000000111110010001011111101011000010111111011101111;//hb2c01f22fd617eef;
		pk[110] = 64'b1101011010010101001011111101100100100100001101101000010100111010;//hd6952fd92436853a;
		pk[111] = 64'b1001000010101100010001111110110010110010011110000101111000000110;//h90ac47ecb2785e06;
		pk[112] = 64'b1001111011001001001001110110101111000000110111001100000100100011;//h9ec9276bc0dcc123;
		pk[113] = 64'b1001000101001011111101100110011111111110101101010100100101100000;//h914bf667feb54960;
		pk[114] = 64'b1010100110101101000110000101110001110110010000011110011100110000;//ha9ad185c7641e730;
		pk[115] = 64'b0111010001011100111010110100101001101111001010011111011110111110;//h745ceb4a6f29f7be;
		pk[116] = 64'b001011010110101110110010110110101001010011000001100101011110;//h2d6bb2da94c195e;
		pk[117] = 64'b1110011011101000111100010000110011000110001101101111010011110000;//he6e8f10cc636f4f0;
		pk[118] = 64'b1010000011001011100111111100110101011110111110010000000100101101;//ha0cb9fcd5ef9012d;
		pk[119] = 64'b0011100101111110101111111100000110110101001111000110111101001111;//h397ebfc1b53c6f4f;
		pk[120] = 64'b0101111010111110011001101010011110100111000000001000100000000111;//h5ebe66a7a7008807;
		pk[121] = 64'b1000001100111001100111101110001011111100110100110100101000100100;//h83399ee2fcd34a24;
		pk[122] = 64'b0111110011110010101010111010101011001001100000101111111010011100;//h7cf2abaac982fe9c;
		pk[123] = 64'b1000_1111_1001_0011_0010_1101_0101_0110_0101_0011_1100_0110_0010_1111_1100_1111;//h8f932d5653c62fcf;

        hash_pk[0] = 64'b1110100110010111110011101011111001110011000101000111100110111010;//'he997cebe731479ba;
        hash_pk[1] = 64'b0001100001111011001110011000011111100110100010111111000110101100;//h187b3987e68bf1ac;
        hash_pk[2] = 64'b0101010111110011100101110100111010101010010010110111011001100000;//h55f3974eaa4b7660;
        hash_pk[3] = 64'b1100001100111010000000001100101011001000111100001010011111011111;//hc33a00cac8f0a7df;

		pseudo_random[0] = 64'b1100010000010000010111110100001111110101000001001111000010110010;//hc4105f43f504f0b2;
		pseudo_random[1] = 64'b1001101111111101011110100100010001001000000100010100010111001101;//h9bfd7a44481145cd;
		pseudo_random[2] = 64'b0011101011010000111000000000110101110111000010011011001010011001;//h3ad0e00d7709b299;
		pseudo_random[3] = 64'b1000110001101000011100011110010101101011101111001011011111001101;//h8c6871e56bbcb7cd;

		ct[0] = 64'b1001001111101111001010011011111101001011001010110101110101001101;//h93ef29bf4b2b5d4d;
		ct[1] = 64'b0111110001110110010001110000111100110000000101110100001101100010;//h7c76470f30174362;
		ct[2] = 64'b0110001111001101000111001111000000001010001010101010100010100011;//h63cd1cf00a2aa8a3;
		ct[3] = 64'b1110111000110001111011110010100101100100010000000101011111110010;//hee31ef29644057f2;
		ct[4] = 64'b1000010010111011000010110111011000010011011001110110101100111001;//h84bb0b7613676b39;
		ct[5] = 64'b0001000010010000110001100100000010101001010001000000010110110100;//h1090c640a94405b4;
		ct[6] = 64'b1111101011000000001100100000110100000111110001100001000110101101;//hfac0320d07c611ad;
		ct[7] = 64'b1111001101010001000011011100010101100000101111000010101010001101;//hf3510dc560bc2a8d;
		ct[8] = 64'b1100111101100000111100100101010000001001110001010000011011100110;//hcf60f25409c506e6;
		ct[9] = 64'b0111010101000011110101111001011100011101111111010000101110111011;//h7543d7971dfd0bbb;
		ct[10] = 64'b1111110001000010100110110000010101111110101110000010011011100110;//hfc429b057eb826e6;
		ct[11] = 64'b0111000000100000101000000001111000001000111000101011111011011111;//h7020a01e08e2bedf;
		ct[12] = 64'b010111001010111010000111011000001101110011100110001100111011;//h5cae8760dce633b;
		ct[13] = 64'b1111111010110100100100101101101110100000110110110001100100100111;//hfeb492dba0db1927;
		ct[14] = 64'b0001111101111010100001010110001010111010101010111001000001011001;//h1f7a8562baab9059;
		ct[15] = 64'b1011001000010010111110100110001111111111011000110001100110101010;//hb212fa63ff6319aa;
		ct[16] = 64'b1000000000101100110001011111001000010000011100100011111100111111;//h802cc5f210723f3f;
		ct[17] = 64'b0010001100111111011101001101011001000011000010010101000000101001;//h233f74d643095029;
		ct[18] = 64'b001111111000100111001001100011100011110101111000011100110001;//h3f89c98e3d78731;
		ct[19] = 64'b1111010101010110010100100011101111110100110100111000011000101111;//hf556523bf4d3862f;
		ct[20] = 64'b0101111001000101001001110000100011000000101110100101000011000010;//h5e452708c0ba50c2;
		ct[21] = 64'b0001101001011111110001110000010111011101111101110101010011011000;//h1a5fc705ddf754d8;
		ct[22] = 64'b1110001001110110000111110001110001010111001111111011001101111100;//he2761f1c573fb37c;
		ct[23] = 64'b1011110111100100000011001110011100010010111110010100110000001101;//hbde40ce712f94c0d;
		ct[24] = 64'b0001000101100001110111011110101001001000100101000111010101001010;//h1161ddea4894754a;
		ct[25] = 64'b1110101110100101001111001000101100001111001001111111111010011011;//heba53c8b0f27fe9b;
		ct[26] = 64'b1110100001000100000111111111110010000000010101000100101010000000;//he8441ffc80544a80;
		ct[27] = 64'b0110111010111000101110100111011001101101111100100000000101001011;//h6eb8ba766df2014b;
		ct[28] = 64'b1111010111110010100010100110010110101110111010110111010111111111;//hf5f28a65aeeb75ff;
		ct[29] = 64'b1011001000110001111100110101101001100010001111101000110010001010;//hb231f35a623e8c8a;
		ct[30] = 64'b1110101100100001011000111010111101100101010111110011010000111001;//heb2163af655f3439;
		ct[31] = 64'b0110100101001110111000000111101000011000110111000100010111001101;//h694ee07a18dc45cd;
		ct[32] = 64'b1100011011010000000111000110110000000010100010000111001010101011;//hc6d01c6c028872ab;
		ct[33] = 64'b0111011100000000011000101011011000110011100100010011011110000110;//h770062b633913786;
		ct[34] = 64'b001101010001100001001001110011111000010110010101110011001001;//h351849cf8595cc9;
		ct[35] = 64'b1100000010010010110111000011001000101101001011000101000101010011;//hc092dc322d2c5153;
		ct[36] = 64'b0101011101001100111000101011011011010100010101100001001000010100;//h574ce2b6d4561214;
		ct[37] = 64'b0101001011100101010101110110011010000110101111111100001001000100;//h52e5576686bfc244;
		ct[38] = 64'b0100010011000110110011100011001100000110011110101111010100001001;//h44c6ce33067af509;
		ct[39] = 64'b1100010001010100111111101010100110010001000011111011110100111110;//hc454fea9910fbd3e;
		ct[40] = 64'b1110000101000000111101001100111110010111100110110001101001000011;//he140f4cf979b1a43;
		ct[41] = 64'b1101011011001011111000001011001110110000010011110000011101111101;//hd6cbe0b3b04f077d;
		ct[42] = 64'b0100101110000101000101111000110101010000101101000000010001000111;//h4b85178d50b40447;
		ct[43] = 64'b0010110001011111010110110111010001110000101011111001000100111010;//h2c5f5b7470af913a;
		ct[44] = 64'b1101110100001100010000100001100101011001011010001010101100001010;//hdd0c42195968ab0a;
		ct[45] = 64'b1101100101110101101011100001010011010100011000000100100001010000;//hd975ae14d4604850;
		ct[46] = 64'b1010100100100100100000111001111000001110100111011101001000011111;//ha924839e0e9dd21f;
		ct[47] = 64'b0001110001111101001011001100101110001011010001001110000111010000;//h1c7d2ccb8b44e1d0;
		ct[48] = 64'b1101100001011000100101000010010111000111011011010001001000100101;//hd8589425c76d1225;
		ct[49] = 64'b0110101000010111101101110010010111001010001010100101001011110000;//h6a17b725ca2a52f0;
		ct[50] = 64'b0101010101100011111110100110001101100110001110001011010100010101;//h5563fa636638b515;
		ct[51] = 64'b0110101111100100011101010011011010001100111011011000000110001001;//h6be475368ced8189;
		ct[52] = 64'b1101000101010111010101110000010011001000001001110001011110000101;//hd1575704c8271785;
		ct[53] = 64'b0100011010000011010001110001100000011110001010100011110100100101;//h468347181e2a3d25;
		ct[54] = 64'b0100110111100011000010110100110001000110010010010110001001110010;//h4de30b4c46496272;
		ct[55] = 64'b1011010000101100010100110111011001011101100110000001010110100111;//hb42c53765d9815a7;
		ct[56] = 64'b100011111000110101101011001110100010101110011101010011000111;    //h8f8d6b3a2b9d4c7;
		ct[57] = 64'b1110101110101000011111101001100100101000011100000101010001101011;//heba87e992870546b;
		ct[58] = 64'b0101000011011001101110000010111001010011100010111110010001111110;//h50d9b82e538be47e;
		ct[59] = 64'b1111000011011000110100110001010100000100111010001110001101111011;//hf0d8d31504e8e37b;
		ct[60] = 64'b0011100111111010010101101110111000110100101111111000101100101011;//h39fa56ee34bf8b2b;
		ct[61] = 64'b1011011100000000001010111101010101111110000011100001101110011111;//hb7002bd57e0e1b9f;
		ct[62] = 64'b0011000110100011110100001110010000010011100110000110101111110110;//h31a3d0e413986bf6;
		ct[63] = 64'b1100000010010101000100010100000100011101011100111000101010011000;//hc09511411d738a98;
		ct[64] = 64'b1100101000110101010011011001111001010010000011101001011100010001;//hca354d9e520e9711;
		ct[65] = 64'b010100001010100000101011011001010000001101100001010010000110;    //h50a82b650361486;
		ct[66] = 64'b011001000011000111100111001011100110000001101101011010100011;    //h6431e72e606d6a3;
		ct[67] = 64'b1100100100100111010000110100000000001101011001000101100100100111;//hc92743400d645927;
		ct[68] = 64'b0110110010001101100101011111110101100110100111110101101100101000;//h6c8d95fd669f5b28;
		ct[69] = 64'b0011011000100001000101011111010010011011010001000011100110101101;//h362115f49b4439ad;
		ct[70] = 64'b0110000101010010011011011101100000100101110001011011111001000100;//h61526dd825c5be44;
		ct[71] = 64'b1110011100101101101100111000010000101011110100011101000111110010;//he72db3842bd1d1f2;
		ct[72] = 64'b110010100010000011110111010110001101111100001010000000111001;//hca20f758df0a039;
		ct[73] = 64'b1011001000001110000010010100100100000111010010101111100011010001;//hb20e0949074af8d1;
		ct[74] = 64'b0001110011001101110101011111100001100010100101011001111110100111;//h1ccdd5f862959fa7;
		ct[75] = 64'b1111011011101001100110000001111000111100000100010100100011000110;//hf6e9981e3c1148c6;
		ct[76] = 64'b0100101101111011110001011100010111011110001011010100001100100110;//h4b7bc5c5de2d4326;
		ct[77] = 64'b1011100101010100111001111101011101110001111101111111111100010111;//hb954e7d771f7ff17;
		ct[78] = 64'b0010100000001011011100001011100000001011100011110001100010110000;//h280b70b80b8f18b0;
		ct[79] = 64'b1100000011100100101110001010101011001011000111011001011111001100;//hc0e4b8aacb1d97cc;
		ct[80] = 64'b0011000000011000100101111110111010001100001001001111010001010110;//h301897ee8c24f456;
		ct[81] = 64'b1110101111100010011001101101011100110001100001010111101100110101;//hebe266d731857b35;
		ct[82] = 64'b0001110100100100101011000111100000110011010010011000110110010101;//h1d24ac7833498d95;
		ct[83] = 64'b1011011101100111010011100000010111001000000010110001001000000101;//hb7674e05c80b1205;
		ct[84] = 64'b0010100011010111011110001000001100010110110110001010010001010000;//h28d7788316d8a450;
		ct[85] = 64'b1010000111110100111101000001011011001011011101001101011000011110;//ha1f4f416cb74d61e;
		ct[86] = 64'b1110101011110010100111110000010000111100010111010101101010110100;//heaf29f043c5d5ab4;
		ct[87] = 64'b0111110001110001010111000001111101001001010010100101101101010010;//h7c715c1f494a5b52;
		ct[88] = 64'b1100110000110001001101100111011101000000011000000100110000010001;//hcc31367740604c11;
		ct[89] = 64'b0101100001000111001011010010001100010000010101000010100101010101;//h58472d2310542955;
		ct[90] = 64'b0001000110011010011001101111001111110110010110100111010010001101;//h119a66f3f65a748d;
		ct[91] = 64'b0001001000010100010110101100010111000111001100011110111011101001;//h12145ac5c731eee9;
		ct[92] = 64'b0101100111110010110111110111110100101000001111010101101000110000;//h59f2df7d283d5a30;
		ct[93] = 64'b1000100100100110100010110000111110000110010110101010011100011101;//h89268b0f865aa71d;
		ct[94] = 64'b1101101111010111111011010111001010000111100110011011110100111011;//hdbd7ed728799bd3b;
		ct[95] = 64'b1100011001011100010010111101100000001011111101000001001101010111;//hc65c4bd80bf41357;
		ct[96] = 64'b101101011011111001001100111110000010110010001111101000011011;//hb5be4cf82c8fa1b;
		ct[97] = 64'b1101111101000111100000100101000100011101011011111100001110111000;//hdf4782511d6fc3b8;
		ct[98] = 64'b0111111001011110100110111101110010011011101001100110110001110010;//h7e5e9bdc9ba66c72;
		ct[99] = 64'b0111001011000000111000111001011101111001010000001100110010011100;//h72c0e3977940cc9c;
		ct[100] = 64'b0111000010001011111001111110110011011010000000111010011110000111;//h708be7ecda03a787;
		ct[101] = 64'b0101100110111010001111101100101001010111001010011011010000100010;//h59ba3eca5729b422;
		ct[102] = 64'b1011110011010000000111100100010001101100100011111100111100011001;//hbcd01e446c8fcf19;
		ct[103] = 64'b0001111111100111011101111101110001110101101101000100111101010111;//h1fe777dc75b44f57;
		ct[104] = 64'b0101111111111011000101001100011010011000000010110110100100111110;//h5ffb14c6980b693e;
		ct[105] = 64'b1010001111001011010111110000000011101011101111110001010101001001;//ha3cb5f00ebbf1549;
		ct[106] = 64'b1010010010010101010001001100100111100001100000001011011010111010;//ha49544c9e180b6ba;
		ct[107] = 64'b0110110010000111110001000000000000010101101010111101000110111000;//h6c87c40015abd1b8;
		ct[108] = 64'b0011110001101001010111101011100001111000001011000011001000011001;//h3c695eb8782c3219;
		ct[109] = 64'b0001011011110010111000110100110111110011011011011001011100110110;//h16f2e34df36d9736;
		ct[110] = 64'b0101001011111010111100111011111010101000110100010000111011101100;//h52faf3bea8d10eec;
		ct[111] = 64'b011000110100000010010100011000111001010111111010110001010111;//h6340946395fac57;
		ct[112] = 64'b1010001000011010011101010111110010101110101111111100010011101110;//ha21a757caebfc4ee;
		ct[113] = 64'b101100001111100011110111101100110010000000110010010100100001;//hb0f8f7b32032521;
		ct[114] = 64'b0100101000010100000110010011110110110111101100110010011110001011;//h4a14193db7b3278b;
		ct[115] = 64'b1000110101100111010110010100110100101000110110100010000101111100;//h8d67594d28da217c;
		ct[116] = 64'b1001111110010011010000110101101100000110000101010111000111001101;//h9f93435b061571cd;
		ct[117] = 64'b0001000001011001100010001110010100010110010001111101110111111101;//h105988e51647ddfd;
		ct[118] = 64'b1101110000101000010100000001110110100011001100000010011011000110;//hdc28501da33026c6;
		ct[119] = 64'b1100100111111111110101111011100010110101001101001101111000000100;//hc9ffd7b8b534de04;
		ct[120] = 64'b1101000011111101101100001111111000011000000100100000010000000101;//hd0fdb0fe18120405;
		ct[121] = 64'b1111100001000101001000001110011010010000010100010010001101001100;//hf84520e69051234c;
		ct[122] = 64'b1110111010100100000110101101010100100001001011101110111101110010;//heea41ad5212eef72;
		ct[123] = 64'b0001110101100011111011101110000010000010110100011010110110001111;//h1d63eee082d1ad8f;
		ct[124] = 64'b1111101000001010111010010000011101010100010100110101111000010011;//hfa0ae90754535e13;
		ct[125] = 64'b1011111110100011111001000011011010010010111101100010010000110010;//hbfa3e43692f62432;
		ct[126] = 64'b1101100010100010000111010101000010011111100110100010001111101110;//hd8a21d509f9a23ee;
		ct[127] = 64'b0101001011001110111011100010000111111101000001111000010100000111;//h52ceee21fd078507;
		ct[128] = 64'b1101100111110001010000000100011011100110101101000100111101011110;//hd9f14046e6b44f5e;
		ct[129] = 64'b1000101101000001011000001001001100100110001111001101110110010101;//h8b416093263cdd95;
		ct[130] = 64'b1000110100110000011001100110010110010010111011101000100011111111;//h8d30666592ee88ff;
		ct[131] = 64'b1101001000110001011101111011011100011101111010100101010111111010;//hd23177b71dea55fa;
		ct[132] = 64'b0010100111001000011110101000110010011011101100100101010011101011;//h29c87a8c9bb254eb;
		ct[133] = 64'b1100000000001101110001010010011111101001001011110100101001011110;//hc00dc527e92f4a5e;
		ct[134] = 64'b1100011100001001010111101110100000101101101001101101110110111011;//hc7095ee82da6ddbb;
		ct[135] = 64'b110000011001011111100010110101100010101111100001110000111010;//hc197e2d62be1c3a;
		
		last_data_on_last_memory_address = 64'b110101;//h35; (in decimal it equals to 53)
		
		set_memory       = 64'b0000000000000000000000000000000000000000000000000000000000000000;



		/// Wait 100 ns for global reset to finish
		#10000000;
        rst = 0;
        
        @(posedge clk1)
        count = 10'd0;
        
        @(posedge clk1)
        crypto_op_1 = 1; crypto_op_2 = 1; crypto_op_3 = 1; // 111 means Execute KEM_DECAPS

/* ------------------------------------------------------------------------------------------------
-- initialize with all memory contents to 0
--------------------------------------------------------------------------------------------------*/      
        
        // Load a 64-bit of 0's to initialize memory contents on all addresses
		for(i=0; i<1024; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = set_memory[j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0; count = i;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            we = 0; addr_ready = 0;
            
            $display("i=%d\n", i);
        end    
        
        $display("starting random seed now");
        
        @(negedge clk1)
        count = 10'd0;

/* ------------------------------------------------------------------------------------------------
-- LOAD pk[i] at memory location [0-123]
--------------------------------------------------------------------------------------------------*/		

        // Load a 64-bit pk[i]
		for(i=0; i<124; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = pk[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end 		

/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Load pseudo_random from 0 to 3 on memory locations #124 to #127
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/	
	
        @(negedge clk1)        
		count = 10'd124;
		
		// Load a 64-bit pseudo_random[i]
		for(i=0; i<4; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = pseudo_random[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end

/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% First 10 values of cpa_secret[i] in memory from #128 to #175
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
        
        @(negedge clk1)        
		count = 10'd128;
		
		// Load a 64-bit cpa_secret[i]
		for(i=0; i<48; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = cpa_secret[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end
        
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Load ct[i] in memory from #200 to #335
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
        
        @(negedge clk1)        
		count = 10'd200;
		
		// Load a 64-bit ct[i]
		for(i=0; i<136; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = ct[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end
        
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Load hash_pk[i] in memory #340-#343
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
        
        @(negedge clk1)        
		count = 10'd340;
		
		// Load a 64-bit hash_pk[i]
		for(i=0; i<4; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = hash_pk[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end
        
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Load a timing counter value at #1023
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/

        // Load a 64-bit timing counter value in memory on #1023 
		for(i=0; i<64; i=i+1)
		begin
			LAD1 = 0; LAD2 = 1;
			@(negedge clk1) 
			din = last_data_on_last_memory_address[i];
		end
		
		@(negedge clk1)
            LAD1 = 0; LAD2 = 0;
		
		// Load a 10-bit corresponding address
		for(i=0; i<10; i=i+1)
		begin
			LAD1 = 1; LAD2 = 0;
			@(negedge clk1) 
			addr = count[i];
		end
		
		// Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
		@(negedge clk1)
		LAD1 = 0; LAD2 = 0;
		
		@(negedge clk1)
		@(negedge clk1)
            we = 1;
            addr_ready = 1;
            
		@(negedge clk1)
		we = 0; addr_ready = 0;
		
/* ------------------------------------------------------------------------------------------------
-- LOAD values ends here
--------------------------------------------------------------------------------------------------*/	
		
		
		/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
		%% Test case to run corresponding operation (i.e. KeyGen, Encaps & Decaps) at once 
		%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
		@(negedge clk1)
		start = 1;	
		@(negedge clk1)
		wait(done);		
		@(negedge clk1)
		start = 0;
		
		/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
		%% Test case to run continuous operation (KeyGen, Encaps, Decaps)
		%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
		
//		@(negedge clk1)
//		start = 1;
//		CONT = 1;
//		#100000;
//		@(negedge clk1)
//		start = 0;
//		$finish();

/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Receiving data onto the chip port as an output
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
	        
        for(count=10'd1008; count<1012; count=count+1)
		begin
                        
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            @(negedge clk1)
                addr_ready = 1;
                    
            for(i=0; i<=66; i=i+1)
            begin
                LAD1 = 1; LAD2 = 1;
                @(negedge clk1);
            end
			
			@(negedge clk1)
                LAD1 = 0; LAD2 = 0;    
        end
        
        $finish();
		
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%%      Test vectors end here for the Decapsulation
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/	       
	end
   
   always #2000  clk1 = ~clk1; 
   always #1000 clk2 = ~clk2; 
      
endmodule
