`timescale 1ns / 1ps

/************************************************************************************************
    1. Design Name:             tb_kem_enc_new
    2. Preparation Date:        June 02, 2021
    3. Initial designed by:     Malik Imran and Samuel Pagliarini (Tallinn University of Technology, Estonia)              
    
    Note! The codes are for academic research use only and does not come with any support or any responsibility. 
****************************************************************************************************/

module tb_kem_enc_new;

	// Inputs to the core
	reg clk1;
	reg clk2;
	reg rst;
	reg addr;
	reg din;
	reg addr_ready;
	reg LAD1;
	reg LAD2;
	reg we;
    reg CONT;
    reg start;	
    reg crypto_op_1;
    reg crypto_op_2;
    reg crypto_op_3;
    	
	// Outputs from the core
	wire dout;
	wire done;
    
	// Registers declaration to hold the test values and signals (i.e., i and count) to drive loops (i.e., for) to read values
	reg [10:0] i;
	reg [9:0] j, count;
	reg [63:0] set_memory;
	reg [63:0] random_seed[3:0];
	reg [63:0] pk[123:0];	// 992 byte pk for SABER_k=3
	
	// Instantiate the Unit Under Test (UUT)	
	wrapper_top uut (
		.clk1(clk1),
		.clk2(clk2), 
		.rst(rst),
		.addr(addr), 
		.din(din), 
		.addr_ready(addr_ready),
		.LAD1(LAD1),
	    .LAD2(LAD2),
	    .we(we),
	    .CONT(CONT),
	    .start(start),
	    .crypto_op_1(crypto_op_1),
	    .crypto_op_2(crypto_op_2), 
	    .crypto_op_3(crypto_op_3),
		.dout(dout),
		.done(done)     		
	);

	initial begin
		// Initialize Inputs
		clk1 = 0;
		clk2 = 0;
		rst = 1;
		addr = 0;
		din = 0;
		addr_ready = 0;
		LAD1 = 0;
		LAD2 = 0;
		we = 0;
		CONT = 0;
		start = 0;
		crypto_op_1 = 0;
	    crypto_op_2 = 0;
	    crypto_op_3 = 0;
	    
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%%      Test vectors for the Encapsulation 
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/	

	
		// 120+4 word pk 
		pk[0] = 64'b1101101100001100101101100111101000010111101010011010111011101011;//hdb0cb67a17a9aeeb;
		pk[1] = 64'b1010111100011001100111111001011011011111101101101110010100100001;//haf199f96dfb6e521;
		pk[2] = 64'b1010100001001100000010110000010110100011000111110000011101110011;//ha84c0b05a31f0773;
		pk[3] = 64'b1110010011100111010110100011100011111110100110110111111010010000;//he4e75a38fe9b7e90;
		pk[4] = 64'b1000001100000110001110111011111101001010101101101111000111101001;//h83063bbf4ab6f1e9;
		pk[5] = 64'b1100111000100100101001111101001101000110000100101001110101100001;//hce24a7d346129d61;
		pk[6] = 64'b0101100111011000011000100111011110110101110001001001001100101100;//h59d86277b5c4932c;
		pk[7] = 64'b1010101011101000010000100110100110001001101000101011111001000111;//haae8426989a2be47;
		pk[8] = 64'b1010001001010001101110101111111111110011101100100111101100011110;//ha251bafff3b27b1e;
		pk[9] =  64'b1100011110101000110000110011001110010001011111111101100110010110;//hc7a8c333917fd996;
		pk[10] = 64'b0010010010110101111001011000110111100011000110001111110101001101;//h24b5e58de318fd4d;
		pk[11] = 64'b1000010000000101011010001001000110000101111010000100000100001110;//h8405689185e8410e;
		pk[12] = 64'b0101001010010000110100011001110011011111010111001100011000100100;//h5290d19cdf5cc624;
		pk[13] = 64'b1000010100011111011100101111011101011010100010101111100000000010;//h851f72f75a8af802;
		pk[14] = 64'b0111110110111001001001111111100111110010011101000100000100000110;//h7db927f9f2744106;
		pk[15] = 64'b0001111110100010000111110010011001011111110011101000000101101001;//h1fa21f265fce8169;
		pk[16] = 64'b0010001110110011011110010011101110111011011101001011111011111010;//h23b3793bbb74befa;
		pk[17] = 64'b1000000110100110101001100000010110100111001000100100100010100101;//h81a6a605a72248a5;
		pk[18] = 64'b0101110010011111011110101111001111010001111011101100001001010111;//h5c9f7af3d1eec257;
		pk[19] = 64'b0011010110111010110000010110011110100110110101011010000101101001;//h35bac167a6d5a169;
		pk[20] = 64'b1011101100110111000111111101001011110001011011111011111111010100;//hbb371fd2f16fbfd4;
		pk[21] = 64'b0011101001001011111011101101110101010101100100110000111000001001;//h3a4beedd55930e09;
		pk[22] = 64'b1010011110110000101000010011100011101000110011001010100010000111;//ha7b0a138e8cca887;
		pk[23] = 64'b100010110010010010000100101101010001010001111010011111110110;//h8b2484b5147a7f6;
		pk[24] = 64'b1101110000110010101000011100110010101111011001001101001110011000;//hdc32a1ccaf64d398;
		pk[25] = 64'b0101110100100011001111000000011100010010111110110101001000001111;//h5d233c0712fb520f;
		pk[26] = 64'b0001101100001010000110110011010000000011011110110001111100101000;//h1b0a1b34037b1f28;
		pk[27] = 64'b0100000111010110110101101101110001100100111011101010011000001011;//h41d6d6dc64eea60b;
		pk[28] = 64'b0110101000101010100010000001111001000111100000100011110100111000;//h6a2a881e47823d38;
		pk[29] = 64'b1010010101010111011101010100001010101000100011101001111110010101;//ha5577542a88e9f95;
		pk[30] = 64'b1101010111010100111100000000010101100101111011101111000010100011;//hd5d4f00565eef0a3;
		pk[31] = 64'b1010100111000010111111101011011000011111000001011001100100101100;//ha9c2feb61f05992c;
		pk[32] = 64'b1010100110111000001001100110011110000011011000010111001101001110;//ha9b826678361734e;
		pk[33] = 64'b0101100011010000000110001001110110101000010110001111010000100111;//h58d0189da858f427;
		pk[34] = 64'b0101011111100001000110010010100011111011110000101001111010011111;//h57e11928fbc29e9f;
		pk[35] = 64'b0010100110001100011000100000101111101100011100101001011101101111;//h298c620bec72976f;
		pk[36] = 64'b1011101001101010101000101110110100110101111111000111110111101000;//hba6aa2ed35fc7de8;
		pk[37] = 64'b010110111010011011011100101010101001011001101101010100011101;//h5ba6dcaa966d51d;
		pk[38] = 64'b0101101100100010000010010110010011001111110011011001110001010001;//h5b220964cfcd9c51;
		pk[39] = 64'b0010110100001011110010100100001100111111000101010111011000011000;//h2d0bca433f157618;
		pk[40] = 64'b1001101101000100001110101010010110100101100101111001011011101111;//h9b443aa5a59796ef;
		pk[41] = 64'b0100111000000101001111111011110010100111111010101110000101000110;//h4e053fbca7eae146;
		pk[42] = 64'b1010000001101110000010001000110010110110001110101010100001011101;//ha06e088cb63aa85d;
		pk[43] = 64'b1011010011101001011001010010100100110010100011001010100111001001;//hb4e96529328ca9c9;
		pk[44] = 64'b0010001111000110100000110001101111000110010100100110110101000110;//h23c6831bc6526d46;
		pk[45] = 64'b1100100110110101010011001110000110001011101000101110111001000101;//hc9b54ce18ba2ee45;
		pk[46] = 64'b0111011001100000111011111111011100011110010001110100010101101111;//h7660eff71e47456f;
		pk[47] = 64'b1001100110001000101010001010011100111111110111111110001110101111;//h9988a8a73fdfe3af;
		pk[48] = 64'b1000100011011111101111111101110010111111001100100010111011000110;//h88dfbfdcbf322ec6;
		pk[49] = 64'b1010001000010000100011001000000000010011010001010110010010010111;//ha2108c8013456497;
		pk[50] = 64'b1110011010010100111010101111011100111000111110101011111100001001;//he694eaf738fabf09;
		pk[51] = 64'b1111111110101101101110001100001110011011000100110000111110101100;//hffadb8c39b130fac;
		pk[52] = 64'b0011110110111110001100000101011001110100001101101010111111000100;//h3dbe30567436afc4;
		pk[53] = 64'b1111111010011100100101110111111001110111001110000101000010100111;//hfe9c977e773850a7;
		pk[54] = 64'b1101110000011100000011100100011100011001101111011100010011000000;//hdc1c0e4719bdc4c0;
		pk[55] = 64'b0111000011111011010000101011001011011100100001100010100100101111;//h70fb42b2dc86292f;
		pk[56] = 64'b1011100100001101001110110111010100101110001100110101011001111111;//hb90d3b752e33567f;
		pk[57] = 64'b1111000111000010100001111001011100001000110000010110100010001110;//hf1c2879708c1688e;
		pk[58] = 64'b1000100101010010000111000000001010001110001111111011001111011011;//h89521c028e3fb3db;
		pk[59] = 64'b1110011001001111001001110110000101100101000011010100010011010110;//he64f2761650d44d6;
		pk[60] = 64'b0011101000111001110010011011111100000001100001100001010011111111;//h3a39c9bf018614ff;
		pk[61] = 64'b0111010010100010000100010001101011011111101010010101000000011010;//h74a2111adfa9501a;
		pk[62] = 64'b1100001011101001000100100100100111110000011010111000000001000111;//hc2e91249f06b8047;
		pk[63] = 64'b0100001111001001100011101011101011100111001101010011110000010000;//h43c98ebae7353c10;
		pk[64] = 64'b1001101010011111110101111010000010101110110110101011010000110010;//h9a9fd7a0aedab432;
		pk[65] = 64'b0100011010110001010101110000100101000101011111101010110100100001;//h46b15709457ead21;
		pk[66] = 64'b0100111101011110111001100111011101000111101001000011101110001101;//h4f5ee67747a43b8d;
		pk[67] = 64'b0011101100001101100100001100111010000000000100001011010000110100;//h3b0d90ce8010b434;
		pk[68] = 64'b0100011001010001101000100111000101101001111010110100011011001011;//h4651a27169eb46cb;
		pk[69] = 64'b1100100011100001101011000000110000011101101010010101101110111101;//hc8e1ac0c1da95bbd;
		pk[70] = 64'b0100100111100110101111001111000100010000011000100011101100110000;//h49e6bcf110623b30;
		pk[71] = 64'b1000101011001110011000010001000011101101100100101111110111001100;//h8ace6110ed92fdcc;
		pk[72] = 64'b1110001011011110111001011100100010001001111001101000111101000110;//he2dee5c889e68f46;
		pk[73] = 64'b1011001111000001100010000001101011110111010111000010110110001100;//hb3c1881af75c2d8c;
		pk[74] = 64'b110100101001100101111001101100000011100000100100001011111101;//hd29979b038242fd;
		pk[75] = 64'b0001110011001110111000000000001001011010110111000010001111101001;//h1ccee0025adc23e9;
		pk[76] = 64'b0111101000100010010010110101000001010100101011110110111001101111;//h7a224b5054af6e6f;
		pk[77] = 64'b1111010110011100011110010100101000011001001111000001100001000100;//hf59c794a193c1844;
		pk[78] = 64'b1000100010111011010100100110101001111101000000011111101101110000;//h88bb526a7d01fb70;
		pk[79] = 64'b1101111100010111101100111111110111000000011000101111100011011111;//hdf17b3fdc062f8df;
		pk[80] = 64'b10011001100110100101011101001100001110100101101111011011;//h999a574c3a5bdb;
		pk[81] = 64'b0110101010001010100001111100110110100000000001010100011100100011;//h6a8a87cda0054723;
		pk[82] = 64'b1000111000010101110010110100101100000110111010011111000100100011;//h8e15cb4b06e9f123;
		pk[83] = 64'b1110100100111100010111110111010101101000111001001101011110010010;//he93c5f7568e4d792;
		pk[84] = 64'b0110101111101001100100110000111000100100110110010010110001101101;//h6be9930e24d92c6d;
		pk[85] = 64'b1011011101001011011011110010001101000010011100111100011011101111;//hb74b6f234273c6ef;
		pk[86] = 64'b0110110110010101111100001001001010100101001101010101010011111110;//h6d95f092a53554fe;
		pk[87] = 64'b0110001100001001000111001100001010001001110110010111000011110010;//h63091cc289d970f2;
		pk[88] = 64'b1010110101000010111110111011001011001001010110101100011001011110;//had42fbb2c95ac65e;
		pk[89] = 64'b1111101110101101101010001110001110001001101001001101011010101011;//hfbada8e389a4d6ab;
		pk[90] = 64'b1011101001110010011111101001011001011110110001010011101111110001;//hba727e965ec53bf1;
		pk[91] = 64'b0101111010101101111101010000010010000101110011001100110110100101;//h5eadf50485cccda5;
		pk[92] = 64'b1011110000001100100011110101011011111111110011001000000011100001;//hbc0c8f56ffcc80e1;
		pk[93] = 64'b0100010111011011100100001101001011111110000000100011001111001111;//h45db90d2fe0233cf;
		pk[94] = 64'b1110110001000001110011110110100100010010100000011010110100010001;//hec41cf691281ad11;
		pk[95] = 64'b1111000101010100101100011001001001011011000011101010111010011100;//hf154b1925b0eae9c;
		pk[96] = 64'b1100111100101001111101100100110100111000110100101101010111000110;//hcf29f64d38d2d5c6;
		pk[97] = 64'b1101001100101111011111100101010011000000110110100000000010101010;//hd32f7e54c0da00aa;
		pk[98] = 64'b0011001110100000110101011101011111011010111000111111111001111100;//h33a0d5d7dae3fe7c;
		pk[99] =  64'b1110000001001101010100111010111011001101110011000011011111110110;//he04d53aecdcc37f6;
		pk[100] = 64'b0001011111010110100001110011110100101010100100101110011000001001;//h17d6873d2a92e609;
		pk[101] = 64'b0101111010100101010111001000100001010010010001100110011001110110;//h5ea55c8852466676;
		pk[102] = 64'b1010100101100110111011001010101110111011101010111001101010110011;//ha966ecabbbab9ab3;
		pk[103] = 64'b1100000000111101010111110100100000101101100000100111000111001101;//hc03d5f482d8271cd;
		pk[104] = 64'b0010011010111111001001010101100101101000110111011111011010100000;//h26bf255968ddf6a0;
		pk[105] = 64'b0111110011000000001011001100001001010011100010001110010000110100;//h7cc02cc25388e434;
		pk[106] = 64'b1101101100000111001111011011100101011110001111110001101010110001;//hdb073db95e3f1ab1;
		pk[107] = 64'b1110101011101000000000010011010001100011100101111000010010111001;//heae80134639784b9;
		pk[108] = 64'b001111011000011101110000110000111111101100000000011100010110;//h3d8770c3fb00716;
		pk[109] = 64'b1011001011000000000111110010001011111101011000010111111011101111;//hb2c01f22fd617eef;
		pk[110] = 64'b1101011010010101001011111101100100100100001101101000010100111010;//hd6952fd92436853a;
		pk[111] = 64'b1001000010101100010001111110110010110010011110000101111000000110;//h90ac47ecb2785e06;
		pk[112] = 64'b1001111011001001001001110110101111000000110111001100000100100011;//h9ec9276bc0dcc123;
		pk[113] = 64'b1001000101001011111101100110011111111110101101010100100101100000;//h914bf667feb54960;
		pk[114] = 64'b1010100110101101000110000101110001110110010000011110011100110000;//ha9ad185c7641e730;
		pk[115] = 64'b0111010001011100111010110100101001101111001010011111011110111110;//h745ceb4a6f29f7be;
		pk[116] = 64'b001011010110101110110010110110101001010011000001100101011110;//h2d6bb2da94c195e;
		pk[117] = 64'b1110011011101000111100010000110011000110001101101111010011110000;//he6e8f10cc636f4f0;
		pk[118] = 64'b1010000011001011100111111100110101011110111110010000000100101101;//ha0cb9fcd5ef9012d;
		pk[119] = 64'b0011100101111110101111111100000110110101001111000110111101001111;//h397ebfc1b53c6f4f;
		pk[120] = 64'b0101111010111110011001101010011110100111000000001000100000000111;//h5ebe66a7a7008807;
		pk[121] = 64'b1000001100111001100111101110001011111100110100110100101000100100;//h83399ee2fcd34a24;
		pk[122] = 64'b0111110011110010101010111010101011001001100000101111111010011100;//h7cf2abaac982fe9c;
		pk[123] = 64'b1000111110010011001011010101011001010011110001100010111111001111;//h8f932d5653c62fcf;
		// 4 word random_seed 
		random_seed[0] = 64'b0000101100000001_1010110101000010_1000000001110001_1001011101111000;//hb01ad4280719778;
		random_seed[1] = 64'b1111000011011110_1101110100010011_0101110111101001_1000101111001001;//hf0dedd135de98bc9;
		random_seed[2] = 64'b1100011110101111_0110111101000010_1001010110101011_0011001101100101;//hc7af6f4295ab3365;
		random_seed[3] = 64'b0110001001000101_1011011110101101_1001100111001101_0111011001001001;//h6245b7ad99cd7649;
		
		set_memory       = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		
		
		// Wait 100 ns for global reset to finish
		#10000000;
        rst = 0;
        
        @(posedge clk1)
        count = 10'd0;
        
        @(posedge clk1)
        crypto_op_1 = 0; crypto_op_2 = 1; crypto_op_3 = 1; // 110 means Execute KEM_ENCAPS

/* ------------------------------------------------------------------------------------------------
-- initialize with all memory contents to 0
--------------------------------------------------------------------------------------------------*/      
        
        // Load a 64-bit of 0's to initialize memory contents on all addresses
		for(i=0; i<1024; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = set_memory[j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0; count = i;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            we = 0; addr_ready = 0;
            
            $display("i=%d\n", i);
        end    
        
        $display("starting random seed now");
        
        @(negedge clk1)
        count = 10'd0;
/* ------------------------------------------------------------------------------------------------
-- LOAD pk[i] at memory location [0-123]
--------------------------------------------------------------------------------------------------*/		

        // Load a 64-bit pk[i]
		for(i=0; i<124; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = pk[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end 
        															
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Load random_seed from 0 to 3
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/	
        @(negedge clk1)        
		count = 10'd140;
		
		// Load a 64-bit random_seed[i]
		for(i=0; i<4; i=i+1)
		begin
            for(j=0; j<64; j=j+1)
            begin
                LAD1 = 0; LAD2 = 1;
                @(negedge clk1) 
                din = random_seed[i][j];
            end
            
            @(negedge clk1)
                LAD1 = 0; LAD2 = 0;
            
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            // Now set write_enable signal to store the loaded data onto a RegFile address inside the ComputeCore3 block
            @(negedge clk1)
            LAD1 = 0; LAD2 = 0;
            
            @(negedge clk1)
            @(negedge clk1)
                we = 1;
                addr_ready = 1;
                
            @(negedge clk1)
            count = count+1; we = 0; addr_ready = 0;
        end 
		
/* ------------------------------------------------------------------------------------------------
-- LOAD values ends here
--------------------------------------------------------------------------------------------------*/
		
		
		/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
		%% Test case to run corresponding operation (i.e. KeyGen, Encaps & Decaps) at once 
		%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
		@(negedge clk1)
		start = 1;	
		@(negedge clk1)
		wait(done);		
		@(negedge clk1)
		start = 0;
		
		/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
		%% Test case to run continuous operation (KeyGen, Encaps, Decaps)
		%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
		
//		@(negedge clk1)
//		start = 1;
//		CONT = 1;
//		#100000;
//		@(negedge clk1)
//		start = 0;
//		$finish();

/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%% Receiving data onto the chip port as an output
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/
	        
        for(count=10'd936; count<940; count=count+1)
		begin
                        
            // Load a 10-bit corresponding address
            for(j=0; j<10; j=j+1)
            begin
                LAD1 = 1; LAD2 = 0;
                @(negedge clk1) 
                addr = count[j];
            end
            
            @(negedge clk1)
                addr_ready = 1;
                    
            for(i=0; i<=66; i=i+1)
            begin
                LAD1 = 1; LAD2 = 1;
                @(negedge clk1);
            end
			
			@(negedge clk1)
                LAD1 = 0; LAD2 = 0;    
        end
        
        $finish();
		
/*%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
%%      Test vectors end here for the Encaps 
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%*/	       
	end
   always #2000  clk1 = ~clk1; 
   always #1000 clk2 = ~clk2; 
      
endmodule
        